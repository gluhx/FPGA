module coder(X, Y);
    //объявляем входы
    input [7:0] X;

    //объявляем выходы
    output [2:0] Y;

    assign Y = (X[7]) ? 3'b111 :
               ((X[6]) ? 3'b110 :
               ((X[5]) ? 3'b101 :
               ((X[4]) ? 3'b100 :
               ((X[3]) ? 3'b011 :
               ((X[2]) ? 3'b010 :
               ((X[1]) ? 3'b001 : 3'b000))))));


endmodule // coder